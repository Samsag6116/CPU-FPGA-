----------------------------------------------------------------------------------------------------------------------------------
--	Copyright <2017> EECE8020 Reconfigurable system Principles. All rights reserved.																	
																																												
--	Summary				:  Lab 5 VHDL code - SHIFTER
--								In this code We use 2 input buses and one function select as a inputs in which function select  
--							   gives what type of operation We want to do on the input(arithmetic or logical) and produce the
--								output and according to that set the status flags(zero, overflow,sign and carry out flags).
								
--	Programmer			:  SAGAR PATEL and EMILY ADAMS
								
--	Revision History	:	01/30/2017 <spatel1652> Rev. <1.0 Initial Creation>
--								02/09/2017 <spatel1652> Rev. <2.0 Commenting the code>

----------------------------------------------------------------------------------------------------------------------------------								

-------------------- Library --------------------

library IEEE;
use IEEE.std_logic_1164.All;
use IEEE.numeric_std.ALL;

-------------------- I/O declaration(entity) --------------------

entity SHIFTER is
port(
		input_bus      : in unsigned   (7 downto 0);
		carry_in       : in std_logic;
		fun_select     : in unsigned	(2 downto 0);
		shifter_output : out unsigned	(7 downto 0);
		carry_out		: out std_logic
		);
end SHIFTER;

-------------------------------- Architecture ---------------------------------------

Architecture RTL of SHIFTER is 

signal temp : unsigned (7 downto 0);

begin

process(fun_select) is

begin
	case (fun_select) is
	
	when ("000") => shifter_output <= input_bus;										--	No shift
  							 carry_out <= carry_in;
							 
	when ("001") => shifter_output <= input_bus sll 1;								-- Shift left
							 carry_out <= carry_in;
			
	when ("010") => shifter_output <= input_bus srl 1;								--	shift Right
							 carry_out <= carry_in;
								 
	when ("011") => shifter_output <="00000000";										-- Put Zeros in output	
							 carry_out <= '0';
								 
	when ("100") => carry_out <= input_bus(7);										-- Rotate left with carry
							 temp <= input_bus sll 1;
							 shifter_output <= temp or ("0000000" & carry_in);
								 
	when ("101") => shifter_output <= input_bus rol 1;								-- rotate left
							 carry_out <= carry_in;
			
	when ("110") => shifter_output <= input_bus ror 1;								-- rotate Right
							 carry_out <= carry_in;
								
	when ("111") => carry_out <= input_bus (0);										-- rotate right with carry
							 temp <= input_bus srl 1;
							 shifter_output <= temp or (carry_in & "0000000");
			
	when others => shifter_output <= input_bus;										-- Display input bus
							carry_out <= carry_in; 
								
		
	end case;
end process;

end RTL;
----------------------------------------------- END --------------------------------------------------